module main

pub fn main() {
	println("Hello from main.v! 😎")
}

pub fn add(a int, b int) int {
	return a + b
}

// pub fn testtest() []int {
// 	arr : []int = [3, 6, 9]
// 	return arr
// 	// return [3, 6, 9]
// }
